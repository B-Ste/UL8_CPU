module top (
    input clk
);

register akku(.clk(clk));
    
endmodule